//module top(
//           input logic clk,
//           input logic reset
//           );
           
//           wire reg_we_E, reg_we_M, reg_we_W;
//           wire[4:0] rd_E, rd_M, rd_W;
//           wire alu_src_E;
//           wire mem_to_reg_E, mem_to_reg_M, mem_to_reg_W;
//           wire[6:0] ALU_control_E;
//           wire[2:0] mem_read_type_E, mem_read_type_M;
//           wire[1:0] mem_store_type_E, mem_store_type_M;
//           wire mem_re_E, mem_re_M;
//           wire[4:0] rs1_E, rs2_E;
//           wire[4:0] rd_E;
//           wire[31:0] imm32_final_E;
//           wire[15:0] pc_E;
//           wire[15:0] pc_plus4E, pc_plus4M;
//           wire branch_flag_M;
//           wire branch_E, branch_M;
//           wire[31:0] read_reg1_E;
//           wire[31:0] read_reg2_E;
//           wire[15:0] dest_pc_E;
//           wire[31:0] ALU_out_M;
//           wire[15
           
           
           